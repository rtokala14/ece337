// $Id: $
// File name:   coefficient_loader.sv
// Created:     3/16/2019
// Author:      ZhiFei Chen
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: coefficient loader
module coefficient_loader(
			input wire clk,
			input wire n_reset,
			input wire new_coefficient_set,
			input wire modwait,
			output reg load_coeff,
			output reg [1:0] coefficient_num);

typedef enum bit [3:0]{IDLE, WAIT0, READY0, WAIT1, READY1, WAIT2, READY2, WAIT3, READY3}stateType;
stateType state;
stateType next_state;

always_ff @(posedge clk, negedge n_reset)begin
	if (n_reset == 0) begin
		state <= IDLE;
	end
	else begin
		state <= next_state;
	end
end

always_comb begin
	next_state = state; //prevent latch
	case(state)
		IDLE: begin
			if((modwait == 0) && (new_coefficient_set == 1))begin
				next_state = WAIT0;
			end
			else begin
				next_state = IDLE;
			end
		end
		WAIT0:begin
			if((modwait == 0))begin
				next_state = READY0;
			end
			else begin
				next_state = WAIT0;
			end
		end
		READY0:begin
			if((modwait == 1))begin
				next_state = WAIT1;
			end
			else begin
				next_state = READY0;
			end
		end
		WAIT1:begin
			if((modwait == 0))begin
				next_state = READY1;
			end
			else begin
				next_state = WAIT1;
			end
		end
		READY1:begin
			if((modwait == 1))begin
				next_state = WAIT2;
			end
			else begin
				next_state = READY1;
			end
		end
		WAIT2:begin
			if((modwait == 0))begin
				next_state = READY2;
			end
			else begin
				next_state = WAIT2;
			end
		end
		READY2:begin
			if((modwait == 1))begin
				next_state = WAIT3;
			end
			else begin
				next_state = READY2;
			end
		end
		WAIT3:begin
			if((modwait == 0))begin
				next_state = READY3;
			end
			else begin
				next_state = WAIT3;
			end
		end
		READY3:begin
			if((modwait == 1))begin
				next_state = IDLE;
			end
			else begin
				next_state = READY3;
			end
		end
	endcase
end //always_comb


always_comb begin
	load_coeff = 1'b0;
	coefficient_num = 2'b00; //prevent latch

	case(state)
		WAIT0:begin
			coefficient_num = 2'b00;
			load_coeff = 1'b0;
		end
		READY0:begin
			coefficient_num = 2'b00;
			load_coeff = 1'b1; //after the coeff loaded 
		end
		WAIT1:begin
			coefficient_num = 2'b01;
			load_coeff = 1'b0;
		end
		READY1:begin
			coefficient_num = 2'b01;
			load_coeff = 1'b1;
		end//after the coeff loaded 
		WAIT2:begin
			coefficient_num = 2'b10;
			load_coeff = 1'b0;
		end
		READY2:begin
			coefficient_num = 2'b10;
			load_coeff = 1'b1;//after the coeff loaded 
		end
		WAIT3:begin
			coefficient_num = 2'b11;
			load_coeff = 1'b0;
		end
		READY3:begin
			coefficient_num = 2'b11;
			load_coeff = 1'b1;
		end
	endcase
end//always comb
endmodule
		
			
