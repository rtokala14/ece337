// $Id: $
// File name:   adder_16bit.sv
// Created:     1/25/2019
// Author:      ZhiFei Chen
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: adder_16bit.
`timescale 1ns / 100ps
module adder_16bit
(
	input wire [15:0] a,
	input wire [15:0] b,
	input wire carry_in,
	output wire [15:0] sum,
	output wire overflow
);
	adder_nbit  #(.BIT_WIDTH(16)) sixteenbit (.a(a), .b(b), .carry_in(carry_in), .sum(sum), .overflow(overflow));
	// STUDENT: Fill in the correct port map with parameter override syntax for using your n-bit ripple carry adder design to be an 8-bit ripple carry adder design
      
	always@*
	  begin
		for(int j = 0; j < 16; j++) begin
		   assert ((( a[j] == 1'b0) || (a[j] == 1'b0)) && ((b[j] == 1'b0) || (b[j] == 1'b1)))
		   else $error("Input  'a' or 'b' of component is not a digital logic value");
		  // #(2) assert ((a[j] + b[j] + carry_in[j]) % 2 == sum[j])
		   //else $error("Output is not correct");
		end
	 end  
endmodule
